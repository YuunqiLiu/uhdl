//[UHDL]Content Start [md5:90afb203fc0f7992cfaf2e6093fdbc66]
module Test (
	input  clk  ,
	input  rst_n);

	//Wire define for this module.

	//Wire define for sub module.

	//Wire define for Inout.

	//Wire sub module connect to this module and inter module connect.

	//Wire this module connect to sub module.

	//module inst.
	test_v comp (
		.clk(clk),
		.rst_n(rst_n));

endmodule
//[UHDL]Content End [md5:90afb203fc0f7992cfaf2e6093fdbc66]

