
module test_v (
    input clk,
    input rst_n
);




endmodule