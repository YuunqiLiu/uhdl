


module module1 #(
    parameter integer unsigned DATA_WIDTH = 32
)(
    input [DATA_WIDTH-1:0] din,
    output [DATA_WIDTH-1:0] dout
);


endmodule